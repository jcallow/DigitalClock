module SevenSegmentDisplay (
							INPUT,
							OUTPUT
							)
							
							
